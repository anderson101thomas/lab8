library verilog;
use verilog.vl_types.all;
entity lastTwoDigits_testbench is
end lastTwoDigits_testbench;
